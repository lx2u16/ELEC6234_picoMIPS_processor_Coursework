//-----------------------------------------------------
// File Name : alucodes.sv
// FuncRon : pMIPS ALU funcRon code definiRons
// Author: tjk
// Last rev. 23 Oct 12
//-----------------------------------------------------
//
`define RA 3'b000
`define RB 3'b001
`define RADD 3'b010
`define RSUB 3'b011
`define RAND 3'b100
`define ROR 3'b101
`define RXOR 3'b110
`define RNOR 3'b111