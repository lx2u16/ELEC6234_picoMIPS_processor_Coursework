`define RB   2'b00
`define RADD 2'b01
`define RMUL 2'b10