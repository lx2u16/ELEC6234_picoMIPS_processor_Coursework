`define NOP  3'b000
`define IN   3'b100
`define ADD  3'b001
`define MULI 3'b110
`define ADDI 3'b101